--Thais Cartuche
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY TB_Ejer3_4 IS
END TB_Ejer3_4;
 
ARCHITECTURE behavior OF TB_Ejer3_4 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Ejer3_4
    PORT(
         CLK : IN  std_logic;
         Q : OUT  std_logic_vector(3 downto 0));
    END COMPONENT;
    

   --Inputs
   signal CLK : std_logic := '0';

 	--Outputs
   signal Q : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Ejer3_4 PORT MAP (
          CLK => CLK,
          Q => Q
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      wait for clk_period;
      wait;
   end process;

END;
